* Unit Inverter
.subckt inv supply Inp Output
* This subcircuit defines a CMOS inverter with equal n and p widths 

.param Wp = 1.91U
.param Wn = 0.665U
.param L = 0.18U
MP1 Output Inp Supply Supply cmosp
+ L=L W=Wp AD = (2*L*Wp) AS = (2*L*Wp) PD = (2*(2*L+Wp)) PS = (2*(2*L+Wp))
MN1 Output Inp 0 0 cmosn
+ L=L W=Wn AD = (2*L*Wn) AS = (2*L*Wn) PD = (2*(2*L+Wn)) PS = (2*(2*L+Wn))
.ends

vdd supply 0 dc 1.8

* Device under test
x3 supply Ck dutout inv

* Load Capacitor
C3 dutout 0 0.05pF

.include models-180nm

*TRANSIENT ANALYSIS with pulse inputs
VCk Ck 0 DC 0 PULSE(0 1.8 0nS 20pS 20pS 4nS 8.0nS)
.tran 1pS 35nS 0nS

.control
run

plot 4.0+V(Ck) V(dutout)
meas tran inrise TRIG v(ck) VAL=0.18 RISE=2 TARG v(Ck) VAL=1.62 RISE=2
meas tran infall TRIG v(ck) VAL=1.62 FALL=2 TARG v(Ck) VAL=0.18 FALL=2
meas tran drise TRIG v(dutout) VAL=0.18 RISE=2 TARG v(dutout) VAL=1.62 RISE=2
meas tran dfall TRIG v(dutout) VAL=1.62 FALL=2 TARG v(dutout) VAL=0.18 FALL=2

.endc
.end
